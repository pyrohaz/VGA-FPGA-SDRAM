-- asmi.vhd

-- Generated using ACDS version 15.1 185

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity asmi is
	port (
		asdo_in             : in  std_logic := '0'; --             asdo_in.sdoin
		asmi_access_granted : in  std_logic := '0'; -- asmi_access_granted.asmi_access_granted
		asmi_access_request : out std_logic;        -- asmi_access_request.asmi_access_request
		data0_out           : out std_logic;        --           data0_out.data0out
		dclk_in             : in  std_logic := '0'; --             dclk_in.dclkin
		ncso_in             : in  std_logic := '0'; --             ncso_in.scein
		noe_in              : in  std_logic := '0'  --              noe_in.noe
	);
end entity asmi;

architecture rtl of asmi is
	component altera_serial_flash_loader is
		generic (
			INTENDED_DEVICE_FAMILY  : string  := "";
			ENHANCED_MODE           : boolean := true;
			ENABLE_SHARED_ACCESS    : string  := "OFF";
			ENABLE_QUAD_SPI_SUPPORT : boolean := false;
			NCSO_WIDTH              : integer := 1
		);
		port (
			dclk_in             : in  std_logic := 'X'; -- dclkin
			ncso_in             : in  std_logic := 'X'; -- scein
			asdo_in             : in  std_logic := 'X'; -- sdoin
			noe_in              : in  std_logic := 'X'; -- noe
			asmi_access_granted : in  std_logic := 'X'; -- asmi_access_granted
			data0_out           : out std_logic;        -- data0out
			asmi_access_request : out std_logic         -- asmi_access_request
		);
	end component altera_serial_flash_loader;

begin

	serial_flash_loader_0 : component altera_serial_flash_loader
		generic map (
			INTENDED_DEVICE_FAMILY  => "Cyclone IV E",
			ENHANCED_MODE           => true,
			ENABLE_SHARED_ACCESS    => "ON",
			ENABLE_QUAD_SPI_SUPPORT => false,
			NCSO_WIDTH              => 1
		)
		port map (
			dclk_in             => dclk_in,             --             dclk_in.dclkin
			ncso_in             => ncso_in,             --             ncso_in.scein
			asdo_in             => asdo_in,             --             asdo_in.sdoin
			noe_in              => noe_in,              --              noe_in.noe
			asmi_access_granted => asmi_access_granted, -- asmi_access_granted.asmi_access_granted
			data0_out           => data0_out,           --           data0_out.data0out
			asmi_access_request => asmi_access_request  -- asmi_access_request.asmi_access_request
		);

end architecture rtl; -- of asmi
